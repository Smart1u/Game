    ����          FAssembly-CSharp, Version=0.0.0.0, Culture=neutral, PublicKeyToken=null   Save+Position   xyzxryrzrwrxcammexpexphealth	maxhealthlevelmoney
skillpointarmorvampirskill
speedskillswordparmorpplayerdamagewin                         Q�DB-�'A>>B    3M>    ��z?�>�      d   d                          d   �  
    